module andGate(out, in1, in2);
        
    input [31:0] in1;
    input [31:0] in2;


    output [31:0] out;

    and AND1(out[0], in1[0], in2[0]);
    and AND2(out[1], in1[1], in2[1]);
    and AND3(out[2], in1[2], in2[2]);
    and AND4(out[3], in1[3], in2[3]);
    and AND5(out[4], in1[4], in2[4]);
    and AND6(out[5], in1[5], in2[5]);
    and AND7(out[6], in1[6], in2[6]);
    and AND8(out[7], in1[7], in2[7]);
    and AND9(out[8], in1[8], in2[8]);
    and AND10(out[9], in1[9], in2[9]);
    and AND11(out[10], in1[10], in2[10]);
    and AND12(out[11], in1[11], in2[11]);
    and AND13(out[12], in1[12], in2[12]);
    and AND14(out[13], in1[13], in2[13]);
    and AND15(out[14], in1[14], in2[14]);
    and AND16(out[15], in1[15], in2[15]);
    and AND17(out[16], in1[16], in2[16]);
    and AND18(out[17], in1[17], in2[17]);
    and AND19(out[18], in1[18], in2[18]);
    and AND20(out[19], in1[19], in2[19]);
    and AND21(out[20], in1[20], in2[20]);
    and AND22(out[21], in1[21], in2[21]);
    and AND23(out[22], in1[22], in2[22]);
    and AND24(out[23], in1[23], in2[23]);
    and AND25(out[24], in1[24], in2[24]);
    and AND26(out[25], in1[25], in2[25]);
    and AND27(out[26], in1[26], in2[26]);
    and AND28(out[27], in1[27], in2[27]);
    and AND29(out[28], in1[28], in2[28]);
    and AND30(out[29], in1[29], in2[29]);
    and AND31(out[30], in1[30], in2[30]);
    and AND32(out[31], in1[31], in2[31]);
    
    // add your code here:

endmodule