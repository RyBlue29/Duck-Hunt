module notGate(out, in);
        
    input [31:0] in;
    output [31:0] out;

    not NOT1(out[0], in[0]);
    not NOT2(out[1], in[1]);
    not NOT3(out[2], in[2]);
    not NOT4(out[3], in[3]);
    not NOT5(out[4], in[4]);
    not NOT6(out[5], in[5]);
    not NOT7(out[6], in[6]);
    not NOT8(out[7], in[7]);
    not NOT9(out[8], in[8]);
    not NOT10(out[9], in[9]);
    not NOT11(out[10], in[10]);
    not NOT12(out[11], in[11]);
    not NOT13(out[12], in[12]);
    not NOT14(out[13], in[13]);
    not NOT15(out[14], in[14]);
    not NOT16(out[15], in[15]);
    not NOT17(out[16], in[16]);
    not NOT18(out[17], in[17]);
    not NOT19(out[18], in[18]);
    not NOT20(out[19], in[19]);
    not NOT21(out[20], in[20]);
    not NOT22(out[21], in[21]);
    not NOT23(out[22], in[22]);
    not NOT24(out[23], in[23]);
    not NOT25(out[24], in[24]);
    not NOT26(out[25], in[25]);
    not NOT27(out[26], in[26]);
    not NOT28(out[27], in[27]);
    not NOT29(out[28], in[28]);
    not NOT30(out[29], in[29]);
    not NOT31(out[30], in[30]);
    not NOT32(out[31], in[31]);


endmodule